module testmod

fn init(){
	println("testmod init")
}

pub fn test() int {
		return 3
}