module main

import os

fn main() {
}